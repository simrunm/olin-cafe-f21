module test_mux32;

  logic [4:0] d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15 , d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31;
  logic [4:0] s;
  wire [4:0] y;

  mux32 UUT(.d0(d0), .d1(d1), .d2(d2), .d3(d3), .d4(d4), .d5(d5), .d6(d6), .d7(d7), .d8(d8), .d9(d9), .d10(d10), .d11(d11), .d12(d12), .d13(d13), .d14(d14), .d15(d15), .d16(d16), .d17(d17), .d18(d18), .d19(d19), .d20(d20), .d21(d21), .d22(d22), .d23(23), .d24(d24), .d25(d25), .d26(d26), .d27(d27), .d28(d28), .d29(d29), .d30(d30), .d31(d31), .s(s), .y(y));

  initial begin
    $dumpvars(0, UUT);
    $dumpfile("mux32.vcd");

    $display("d0|d1|d2|d3|d4|d5|d6|d7|d8|d9|d10|d11|d12|d13|d14|d15|d16|d17|d18|d19|d20|d21|d22|d23|d24|d25|d26|d27|d28|d29|d30|d31|s |y");
    // testing three random cases

    for (int i = 0; i < 32; i = i + 1) begin 
      
      d0 = 5'b00000 + i;
      d1 = 5'b00001 + i;
      d2 = 5'b00010 + i;
      d3 = 5'b00011 + i;
      d4 = 5'b00100 + i;
      d5 = 5'b00101 + i;
      d6 = 5'b00110 + i;
      d7 = 5'b00111 + i;
      d8 = 5'b01000 + i;
      d9 = 5'b01001 + i;
      d10 = 5'b01010 + i;
      d11 = 5'b01011 + i;
      d12 = 5'b01100 + i;
      d13 = 5'b01101 + i;
      d14 = 5'b01110 + i;
      d15 = 5'b01111 + i;
      d16 = 5'b10000 + i;
      d17 = 5'b10001 + i;
      d18 = 5'b10010 + i;
      d19 = 5'b10011 + i;
      d20 = 5'b10100 + i;
      d21 = 5'b10101 + i;
      d22 = 5'b10110 + i;
      d23 = 5'b10111 + i;
      d24 = 5'b11000 + i;
      d25 = 5'b11001 + i;
      d26 = 5'b11010 + i;
      d27 = 5'b11011 + i;
      d28 = 5'b11100 + i;
      d29 = 5'b11101 + i;
      d30 = 5'b11110 + i;
      d31 = 5'b11111 + i; 
      s = 5'b00000 + i;
      #1 $display("%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b|%b", d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15 , d16, d17, d18, d19, d20, d21, d22, d23, d24, d25, d26, d27, d28, d29, d30, d31, s, y);
    end
  end

endmodule